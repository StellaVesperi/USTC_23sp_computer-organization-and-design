`timescale 1ns / 1ps

module AND(
input [31:0] lhs, rhs,
output [31:0] res
);
assign res=(lhs&rhs);
endmodule
